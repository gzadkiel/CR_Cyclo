module window_selector_LUT #(
    parameter NP = 1024 //! Number of FFT points parameter
) (
    input   [2         : 0] i_NFFT_sel, //! Input to select number of FFT points
    input   [1         : 0] i_WIND_sel, //! Input to select window type 
    output  [NP*10 - 1 : 0] o_window    //! Packed array with window coefficients
);

always @(*) begin
    // if (i_WIND_sel == NB_SEL'b00) begin // Rectangular
    //     case (i_NFFT_sel)
    //         3'b000 : o_window = {160{1'b1}};
    //         3'b001 : o_window = {320{1'b1}};
    //         3'b010 : o_window = {640{1'b1}};
    //         3'b011 : o_window = {1280{1'b1}};
    //         3'b100 : o_window = {2560{1'b1}};
    //         3'b101 : o_window = {5120{1'b1}};
    //         3'b110 : o_window = {10240{1'b1}}; 
    //     endcase   
    // end
    if (i_WIND_sel == NB_SEL'b01) begin // Hamming
        case (i_NFFT_sel)
            3'b000 : o_window = 160'b0000001010000000111100000111010000110010000100101100011000100001110100000111111000011111100001110100000110001000010010110000110010000001110100000011110000001010;
            3'b001 : o_window = 320'b00000010100000001011000000111100000101000000011100000010010100001100000000111100000100100000010100110001011111000110100100011100010001111000000111110100011111110001111111000111110100011110000001110001000110100100010111110001010011000100100000001111000000110000000010010100000111000000010100000000111100000010110000001010;
            3'b010 : o_window = 640'b0000001010000000101000000010110000001100000000111000000100010000010100000001100000000111000000100000000010010100001010100000101111000011010100001110100001000000000100011000010011000001010010000101011100010111010001100010000110011100011011000001110000000111010000011101110001111010000111110000011111100001111111000111111100011111110001111111000111111000011111000001111010000111011100011101000001110000000110110000011001110001100010000101110100010101110001010010000100110000010001100001000000000011101000001101010000101111000010101000001001010000100000000001110000000110000000010100000001000100000011100000001100000000101100000010100000001010;
            3'b011 : o_window = 1280'b00000010100000001010000000101000000010100000001011000000110000000011000000001101000000111000000011110000010001000001001000000101000000010110000001011100000110010000011011000001110100001000000000100010000010010000001001110000101001000010110000001011110000110001000011010000001101110000111010000011110100010000000001000010000100010100010010000001001011000100111000010100010001010100000101011100010110010001011100000101111100011000010001100100000110011000011010010001101011000110110100011011110001110001000111001100011101010001110110000111100000011110010001111010000111101100011111000001111101000111111000011111110001111111000111111100011111110001111111000111111100011111110001111111000111111000011111010001111100000111101100011110100001111001000111100000011101100001110101000111001100011100010001101111000110110100011010110001101001000110011000011001000001100001000101111100010111000001011001000101011100010101000001010001000100111000010010110001001000000100010100010000100001000000000011110100001110100000110111000011010000001100010000101111000010110000001010010000100111000010010000001000100000100000000001110100000110110000011001000001011100000101100000010100000001001000000100010000001111000000111000000011010000001100000000110000000010110000001010000000101000000010100000001010;
            3'b100 : o_window = 2560'b0000001010000000101000000010100000001010000000101000000010100000001010000000101100000010110000001011000000110000000011000000001100000000110100000011010000001110000000111000000011110000001111000001000000000100010000010001000001001000000100110000010100000001010100000101010000010110000001011100000110000000011001000001101000000110110000011100000001110100000111100000011111000010000100001000100000100011000010010000001001010000100111000010100000001010010000101010000010110000001011010000101110000011000000001100010000110010000011010000001101010000110111000011100000001110010000111011000011110000001111100000111111000100000100010000100001000100000100010100010001100001001000000100100100010010110001001100000100111000010011110001010001000101001000010100110001010101000101011000010110000001011001000101101000010111000001011101000101111000011000000001100001000110001000011000110001100101000110011000011001110001101000000110100100011010100001101011000110110100011011100001101111000111000000011100010001110010000111001000011100110001110100000111010100011101100001110111000111011100011110000001111001000111100100011110100001111011000111101100011111000001111100000111110100011111010001111110000111111000011111100001111110000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111110000111111000011111100001111110000111110100011111010001111100000111110000011110110001111011000111101000011110010001111001000111100000011101110001110111000111011000011101010001110100000111001100011100100001110010000111000100011100000001101111000110111000011011010001101011000110101000011010010001101000000110011100011001100001100101000110001100011000100001100001000110000000010111100001011101000101110000010110100001011001000101100000010101100001010101000101001100010100100001010001000100111100010011100001001100000100101100010010010001001000000100011000010001010001000100000100001000010000010000111111000011111000001111000000111011000011100100001110000000110111000011010100001101000000110010000011000100001100000000101110000010110100001011000000101010000010100100001010000000100111000010010100001001000000100011000010001000001000010000011111000001111000000111010000011100000001101100000110100000011001000001100000000101110000010110000001010100000101010000010100000001001100000100100000010001000001000100000100000000001111000000111100000011100000001110000000110100000011010000001100000000110000000011000000001011000000101100000010110000001010000000101000000010100000001010000000101000000010100000001010;
            3'b101 : o_window = 5120'b00000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101100000010110000001011000000101100000010110000001011000000110000000011000000001100000000110000000011000000001101000000110100000011010000001101000000110100000011100000001110000000111000000011110000001111000000111100000011110000010000000001000000000100000000010001000001000100000100010000010010000001001000000100110000010011000001001100000101000000010100000001010100000101010000010101000001011000000101100000010111000001011100000110000000011000000001100100000110010000011010000001101000000110110000011011000001110000000111000000011101000001110100000111100000011110000001111100000111110000100000000010000000001000010000100010000010001000001000110000100011000010010000001001010000100101000010011000001001100000100111000010100000001010000000101001000010101000001010100000101011000010110000001011000000101101000010111000001011100000101111000011000000001100000000110001000011001000001100100000110011000011010000001101000000110101000011011000001101100000110111000011100000001110010000111001000011101000001110110000111011000011110000001111010000111110000011111000001111110001000000000100000000010000010001000010000100001100010000110001000100000100010100010001100001000110000100011100010010000001001000000100100100010010100001001011000100101100010011000001001101000100110100010011100001001111000101000000010100000001010001000101001000010100100001010011000101010000010101010001010101000101011000010101110001010111000101100000010110010001011001000101101000010110110001011011000101110000010111010001011101000101111000010111110001011111000110000000011000010001100001000110001000011000100001100011000110010000011001000001100101000110011000011001100001100111000110011100011010000001101000000110100100011010100001101010000110101100011010110001101100000110110000011011010001101101000110111000011011100001101111000110111100011100000001110000000111000100011100010001110010000111001000011100110001110011000111010000011101000001110101000111010100011101010001110110000111011000011101110001110111000111011100011110000001111000000111100000011110010001111001000111100100011110100001111010000111101000011110110001111011000111101100011110110001111100000111110000011111000001111100000111110100011111010001111101000111110100011111010001111110000111111000011111100001111110000111111000011111100001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111110000111111000011111100001111110000111111000011111100001111101000111110100011111010001111101000111110100011111000001111100000111110000011111000001111011000111101100011110110001111011000111101000011110100001111010000111100100011110010001111001000111100000011110000001111000000111011100011101110001110111000111011000011101100001110101000111010100011101010001110100000111010000011100110001110011000111001000011100100001110001000111000100011100000001110000000110111100011011110001101110000110111000011011010001101101000110110000011011000001101011000110101100011010100001101010000110100100011010000001101000000110011100011001110001100110000110011000011001010001100100000110010000011000110001100010000110001000011000010001100001000110000000010111110001011111000101111000010111010001011101000101110000010110110001011011000101101000010110010001011001000101100000010101110001010111000101011000010101010001010101000101010000010100110001010010000101001000010100010001010000000101000000010011110001001110000100110100010011010001001100000100101100010010110001001010000100100100010010000001001000000100011100010001100001000110000100010100010001000001000011000100001100010000100001000001000100000000010000000000111111000011111000001111100000111101000011110000001110110000111011000011101000001110010000111001000011100000001101110000110110000011011000001101010000110100000011010000001100110000110010000011001000001100010000110000000011000000001011110000101110000010111000001011010000101100000010110000001010110000101010000010101000001010010000101000000010100000001001110000100110000010011000001001010000100101000010010000001000110000100011000010001000001000100000100001000010000000001000000000011111000001111100000111100000011110000001110100000111010000011100000001110000000110110000011011000001101000000110100000011001000001100100000110000000011000000001011100000101110000010110000001011000000101010000010101000001010100000101000000010100000001001100000100110000010011000001001000000100100000010001000001000100000100010000010000000001000000000100000000001111000000111100000011110000001111000000111000000011100000001110000000110100000011010000001101000000110100000011010000001100000000110000000011000000001100000000110000000010110000001011000000101100000010110000001011000000101100000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010;
            3'b110 : o_window = 10240'b0000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001011000000101100000010110000001011000000101100000010110000001011000000101100000010110000001011000000101100000010110000001011000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001101000000110100000011010000001101000000110100000011010000001101000000110100000011100000001110000000111000000011100000001110000000111000000011100000001111000000111100000011110000001111000000111100000011110000001111000001000000000100000000010000000001000000000100000000010000000001000100000100010000010001000001000100000100010000010001000001001000000100100000010010000001001000000100100000010011000001001100000100110000010011000001001100000100110000010100000001010000000101000000010100000001010100000101010000010101000001010100000101010000010110000001011000000101100000010110000001011000000101110000010111000001011100000101110000011000000001100000000110000000011000000001100100000110010000011001000001100100000110100000011010000001101000000110100000011011000001101100000110110000011011000001110000000111000000011100000001110000000111010000011101000001110100000111010000011110000001111000000111100000011110000001111100000111110000011111000010000000001000000000100000000010000000001000010000100001000010000100001000100000100010000010001000001000100000100011000010001100001000110000100100000010010000001001000000100101000010010100001001010000100101000010011000001001100000100110000010011100001001110000100111000010100000001010000000101000000010100100001010010000101001000010101000001010100000101010000010101100001010110000101011000010110000001011000000101100000010110000001011010000101101000010110100001011100000101110000010111000001011110000101111000010111100001100000000110000000011000100001100010000110001000011001000001100100000110010000011001100001100110000110011000011010000001101000000110100000011010100001101010000110101000011011000001101100000110110000011011100001101110000110111000011100000001110000000111001000011100100001110010000111010000011101000001110100000111011000011101100001110110000111100000011110000001111000000111101000011110100001111010000111110000011111000001111110000111111000011111100010000000001000000000100000000010000010001000001000100000100010000100001000010000100001100010000110001000011000100010000010001000001000100000100010100010001010001000101000100011000010001100001000111000100011100010001110001001000000100100000010010000001001001000100100100010010010001001010000100101000010010100001001011000100101100010011000001001100000100110000010011010001001101000100110100010011100001001110000100111000010011110001001111000100111100010100000001010000000101000100010100010001010001000101001000010100100001010010000101001100010100110001010011000101010000010101000001010100000101010100010101010001010101000101011000010101100001010111000101011100010101110001011000000101100000010110000001011001000101100100010110010001011010000101101000010110100001011011000101101100010110110001011100000101110000010111000001011101000101110100010111010001011110000101111000010111100001011111000101111100010111110001100000000110000000011000000001100000000110000100011000010001100001000110001000011000100001100010000110001100011000110001100011000110010000011001000001100100000110010100011001010001100101000110010100011001100001100110000110011000011001110001100111000110011100011010000001101000000110100000011010000001101001000110100100011010010001101010000110101000011010100001101010000110101100011010110001101011000110101100011011000001101100000110110000011011010001101101000110110100011011010001101110000110111000011011100001101110000110111100011011110001101111000110111100011100000001110000000111000000011100000001110001000111000100011100010001110001000111001000011100100001110010000111001000011100100001110011000111001100011100110001110011000111010000011101000001110100000111010000011101000001110101000111010100011101010001110101000111010100011101100001110110000111011000011101100001110110000111011100011101110001110111000111011100011101110001111000000111100000011110000001111000000111100000011110000001111001000111100100011110010001111001000111100100011110010001111010000111101000011110100001111010000111101000011110100001111011000111101100011110110001111011000111101100011110110001111011000111101100011111000001111100000111110000011111000001111100000111110000011111000001111100000111110100011111010001111101000111110100011111010001111101000111110100011111010001111101000111111000011111100001111110000111111000011111100001111110000111111000011111100001111110000111111000011111100001111110000111111000011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111100001111110000111111000011111100001111110000111111000011111100001111110000111111000011111100001111110000111111000011111100001111101000111110100011111010001111101000111110100011111010001111101000111110100011111010001111100000111110000011111000001111100000111110000011111000001111100000111110000011110110001111011000111101100011110110001111011000111101100011110110001111011000111101000011110100001111010000111101000011110100001111010000111100100011110010001111001000111100100011110010001111001000111100000011110000001111000000111100000011110000001111000000111011100011101110001110111000111011100011101110001110110000111011000011101100001110110000111011000011101010001110101000111010100011101010001110101000111010000011101000001110100000111010000011101000001110011000111001100011100110001110011000111001000011100100001110010000111001000011100100001110001000111000100011100010001110001000111000000011100000001110000000111000000011011110001101111000110111100011011110001101110000110111000011011100001101110000110110100011011010001101101000110110100011011000001101100000110110000011010110001101011000110101100011010110001101010000110101000011010100001101010000110100100011010010001101001000110100000011010000001101000000110100000011001110001100111000110011100011001100001100110000110011000011001010001100101000110010100011001010001100100000110010000011001000001100011000110001100011000110001100010000110001000011000100001100001000110000100011000010001100000000110000000011000000001100000000101111100010111110001011111000101111000010111100001011110000101110100010111010001011101000101110000010111000001011100000101101100010110110001011011000101101000010110100001011010000101100100010110010001011001000101100000010110000001011000000101011100010101110001010111000101011000010101100001010101000101010100010101010001010100000101010000010101000001010011000101001100010100110001010010000101001000010100100001010001000101000100010100010001010000000101000000010011110001001111000100111100010011100001001110000100111000010011010001001101000100110100010011000001001100000100110000010010110001001011000100101000010010100001001010000100100100010010010001001001000100100000010010000001001000000100011100010001110001000111000100011000010001100001000101000100010100010001010001000100000100010000010001000001000011000100001100010000110001000010000100001000010000010001000001000100000100010000000001000000000100000000001111110000111111000011111100001111100000111110000011110100001111010000111101000011110000001111000000111100000011101100001110110000111011000011101000001110100000111010000011100100001110010000111001000011100000001110000000110111000011011100001101110000110110000011011000001101100000110101000011010100001101010000110100000011010000001101000000110011000011001100001100110000110010000011001000001100100000110001000011000100001100010000110000000011000000001011110000101111000010111100001011100000101110000010111000001011010000101101000010110100001011000000101100000010110000001011000000101011000010101100001010110000101010000010101000001010100000101001000010100100001010010000101000000010100000001010000000100111000010011100001001110000100110000010011000001001100000100101000010010100001001010000100101000010010000001001000000100100000010001100001000110000100011000010001000001000100000100010000010001000001000010000100001000010000100001000000000100000000010000000001000000000011111000001111100000111110000011110000001111000000111100000011110000001110100000111010000011101000001110100000111000000011100000001110000000111000000011011000001101100000110110000011011000001101000000110100000011010000001101000000110010000011001000001100100000110010000011000000001100000000110000000011000000001011100000101110000010111000001011100000101100000010110000001011000000101100000010110000001010100000101010000010101000001010100000101010000010100000001010000000101000000010100000001001100000100110000010011000001001100000100110000010011000001001000000100100000010010000001001000000100100000010001000001000100000100010000010001000001000100000100010000010000000001000000000100000000010000000001000000000100000000001111000000111100000011110000001111000000111100000011110000001111000000111000000011100000001110000000111000000011100000001110000000111000000011010000001101000000110100000011010000001101000000110100000011010000001101000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001011000000101100000010110000001011000000101100000010110000001011000000101100000010110000001011000000101100000010110000001011000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001010; 
        endcase     
    end
    else if (i_WIND_sel == NB_SEL'b10) begin // Blackman
        case (i_NFFT_sel)
            3'b000 : o_window = 160'b1111111111000000001000000010010000011001000011001000010100000001101100000111110100011111010001101100000101000000001100100000011001000000100100000000101111111111;
            3'b001 : o_window = 320'b11111111110000000000000000001000000001000000001001000000111100000101110000100010000010111000001111000001001011000101101000011001110001110011000111101100011111110001111111000111101100011100110001100111000101101000010010110000111100000010111000001000100000010111000000111100000010010000000100000000001000000000001111111111;
            3'b010 : o_window = 640'b1111111111000000000000000000000000000001000000000100000000110000000100000000011000000010000000001011000000111000000100100000010110000001101100001000010000100110000010110100001100110000111010000100000100010010010001010000000101011100010111100001100101000110101100011100010001110101000111100100011111000001111110000111111100011111110001111110000111110000011110010001110101000111000100011010110001100101000101111000010101110001010000000100100100010000010000111010000011001100001011010000100110000010000100000110110000010110000001001000000011100000001011000000100000000001100000000100000000001100000000010000000001000000000000000000001111111111;
            3'b011 : o_window = 1280'b11111111110000000000000000000000000000000000000000000000000000000000010000000001000000000100000000100000000011000000001100000001000000000101000000011000000001110000001000000000100100000010110000001100000000111000000100000000010010000001010000000101100000011000000001101100000111010000100000000010001100001001100000101001000010110000001011110000110010000011011000001110010000111101000100000000010001000001001000000100101100010011110001010011000101011000010110100001011101000110000000011001000001100111000110101000011011010001101111000111001000011101000001110111000111100000011110100001111100000111110100011111100001111111000111111100011111110001111111000111111100011111110001111110000111110100011111000001111010000111100000011101110001110100000111001000011011110001101101000110101000011001110001100100000110000000010111010001011010000101011000010100110001001111000100101100010010000001000100000100000000001111010000111001000011011000001100100000101111000010110000001010010000100110000010001100001000000000011101000001101100000110000000010110000001010000000100100000010000000000111000000011000000001011000000100100000010000000000111000000011000000001010000000100000000001100000000110000000010000000000100000000010000000001000000000000000000000000000000000000000000000000001111111111;
            3'b100 : o_window = 2560'b1111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000010000000001000000000100000000100000000010000000001000000000110000000011000000001100000001000000000100000000010000000001010000000101000000011000000001100000000111000000011100000010000000001001000000100100000010100000001011000000110000000011000000001101000000111000000011110000010000000001000100000100100000010011000001010000000101010000010110000001011100000110000000011001000001101000000111000000011101000001111000001000000000100001000010001000001001000000100101000010011100001010000000101010000010101100001011010000101111000011000000001100100000110100000011010100001101110000111001000011101100001111000000111110000100000000010000100001000011000100010100010001110001001001000100101100010011010001001110000101000000010100100001010100000101011000010101110001011001000101101100010111000001011110000110000000011000010001100011000110010100011001100001101000000110100100011010110001101100000110111000011011110001110000000111000100011100110001110100000111010100011101100001110111000111100000011110010001111010000111101100011110110001111100000111110100011111010001111110000111111000011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111100001111110000111110100011111010001111100000111101100011110110001111010000111100100011110000001110111000111011000011101010001110100000111001100011100010001110000000110111100011011100001101100000110101100011010010001101000000110011000011001010001100011000110000100011000000001011110000101110000010110110001011001000101011100010101100001010100000101001000010100000001001110000100110100010010110001001001000100011100010001010001000011000100001000010000000000111110000011110000001110110000111001000011011100001101010000110100000011001000001100000000101111000010110100001010110000101010000010100000001001110000100101000010010000001000100000100001000010000000000111100000011101000001110000000110100000011001000001100000000101110000010110000001010100000101000000010011000001001000000100010000010000000000111100000011100000001101000000110000000011000000001011000000101000000010010000001001000000100000000001110000000111000000011000000001100000000101000000010100000001000000000100000000010000000000110000000011000000001100000000100000000010000000001000000000010000000001000000000100000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111;
            3'b101 : o_window = 5120'b11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000100000000010000000001000000000100000000010000000001000000000100000000011000000001100000000110000000011000000001100000000110000000100000000010000000001000000000100000000010000000001010000000101000000010100000001010000000110000000011000000001100000000110000000011100000001110000000111000000011100000010000000001000000000100000000010010000001001000000100100000010100000001010000000101000000010110000001011000000101100000011000000001100000000110100000011010000001101000000111000000011100000001111000000111100000100000000010000000001000100000100010000010001000001001000000100100000010011000001001100000101000000010101000001010100000101100000010110000001011100000101110000011000000001100000000110010000011010000001101000000110110000011100000001110000000111010000011101000001111000000111110000011111000010000000001000010000100010000010001000001000110000100100000010010000001001010000100110000010011100001001110000101000000010100100001010100000101010000010101100001011000000101101000010111000001011100000101111000011000000001100010000110010000011001100001100110000110100000011010100001101100000110111000011100000001110010000111001000011101000001110110000111100000011110100001111100000111111000100000000010000000001000001000100001000010000110001000100000100010100010001100001000111000100100000010010010001001010000100101000010010110001001100000100110100010011100001001111000101000000010100010001010010000101001100010100110001010100000101010100010101100001010111000101100000010110010001011010000101101000010110110001011100000101110100010111100001011111000110000000011000000001100001000110001000011000110001100100000110010000011001010001100110000110011100011010000001101000000110100100011010100001101010000110101100011011000001101101000110110100011011100001101111000110111100011100000001110001000111000100011100100001110010000111001100011101000001110100000111010100011101010001110110000111011000011101110001110111000111100000011110000001111001000111100100011110100001111010000111101000011110110001111011000111110000011111000001111100000111110100011111010001111101000111110100011111100001111110000111111000011111100001111110000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111100001111110000111111000011111100001111110000111110100011111010001111101000111110100011111000001111100000111110000011110110001111011000111101000011110100001111010000111100100011110010001111000000111100000011101110001110111000111011000011101100001110101000111010100011101000001110100000111001100011100100001110010000111000100011100010001110000000110111100011011110001101110000110110100011011010001101100000110101100011010100001101010000110100100011010000001101000000110011100011001100001100101000110010000011001000001100011000110001000011000010001100000000110000000010111110001011110000101110100010111000001011011000101101000010110100001011001000101100000010101110001010110000101010100010101000001010011000101001100010100100001010001000101000000010011110001001110000100110100010011000001001011000100101000010010100001001001000100100000010001110001000110000100010100010001000001000011000100001000010000010001000000000100000000001111110000111110000011110100001111000000111011000011101000001110010000111001000011100000001101110000110110000011010100001101000000110011000011001100001100100000110001000011000000001011110000101110000010111000001011010000101100000010101100001010100000101010000010100100001010000000100111000010011100001001100000100101000010010000001001000000100011000010001000001000100000100001000010000000000111110000011111000001111000000111010000011101000001110000000111000000011011000001101000000110100000011001000001100000000110000000010111000001011100000101100000010110000001010100000101010000010100000001001100000100110000010010000001001000000100010000010001000001000100000100000000010000000000111100000011110000001110000000111000000011010000001101000000110100000011000000001100000000101100000010110000001011000000101000000010100000001010000000100100000010010000001001000000100000000010000000001000000000011100000001110000000111000000011100000001100000000110000000011000000001100000000101000000010100000001010000000101000000010000000001000000000100000000010000000001000000000011000000001100000000110000000011000000001100000000110000000010000000001000000000100000000010000000001000000000100000000010000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111;
            3'b110 : o_window = 10240'b1111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001100000000110000000011000000001100000000110000000011000000001100000000110000000011100000001110000000111000000011100000001110000000111000000011100000010000000001000000000100000000010000000001000000000100000000010000000001001000000100100000010010000001001000000100100000010010000001010000000101000000010100000001010000000101000000010110000001011000000101100000010110000001011000000101100000011000000001100000000110000000011000000001100000000110100000011010000001101000000110100000011010000001110000000111000000011100000001110000000111000000011110000001111000000111100000011110000010000000001000000000100000000010000000001000000000100010000010001000001000100000100010000010010000001001000000100100000010010000001001100000100110000010011000001001100000101000000010100000001010000000101000000010101000001010100000101010000010110000001011000000101100000010110000001011100000101110000010111000001100000000110000000011000000001100000000110010000011001000001100100000110100000011010000001101000000110110000011011000001101100000110110000011100000001110000000111000000011101000001110100000111010000011110000001111000000111100000011111000001111100000111110000100000000010000000001000000000100001000010000100001000010000100010000010001000001000110000100011000010001100001001000000100100000010010000001001010000100101000010010100001001100000100110000010011100001001110000100111000010100000001010000000101000000010100100001010010000101010000010101000001010100000101011000010101100001011000000101100000010110000001011010000101101000010111000001011100000101110000010111100001011110000110000000011000000001100000000110001000011000100001100100000110010000011001000001100110000110011000011010000001101000000110101000011010100001101010000110110000011011000001101110000110111000011100000001110000000111000000011100100001110010000111010000011101000001110110000111011000011101100001111000000111100000011110100001111010000111110000011111000001111110000111111000011111100010000000001000000000100000100010000010001000010000100001000010000110001000011000100001100010001000001000100000100010100010001010001000110000100011000010001110001000111000100100000010010000001001000000100100100010010010001001010000100101000010010110001001011000100110000010011000001001101000100110100010011010001001110000100111000010011110001001111000101000000010100000001010001000101000100010100010001010010000101001000010100110001010011000101010000010101000001010101000101010100010101010001010110000101011000010101110001010111000101100000010110000001011001000101100100010110010001011010000101101000010110110001011011000101110000010111000001011100000101110100010111010001011110000101111000010111110001011111000101111100011000000001100000000110000100011000010001100001000110001000011000100001100011000110001100011000110001100100000110010000011001010001100101000110010100011001100001100110000110011100011001110001100111000110100000011010000001101001000110100100011010010001101010000110101000011010100001101011000110101100011010110001101100000110110000011011000001101101000110110100011011100001101110000110111000011011110001101111000110111100011100000001110000000111000000011100000001110001000111000100011100010001110010000111001000011100100001110011000111001100011100110001110100000111010000011101000001110100000111010100011101010001110101000111010100011101100001110110000111011000011101110001110111000111011100011101110001110111000111100000011110000001111000000111100000011110010001111001000111100100011110010001111010000111101000011110100001111010000111101000011110110001111011000111101100011110110001111011000111101100011111000001111100000111110000011111000001111100000111110000011111010001111101000111110100011111010001111101000111110100011111010001111110000111111000011111100001111110000111111000011111100001111110000111111000011111100001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111000011111100001111110000111111000011111100001111110000111111000011111100001111110000111110100011111010001111101000111110100011111010001111101000111110100011111000001111100000111110000011111000001111100000111110000011110110001111011000111101100011110110001111011000111101100011110100001111010000111101000011110100001111010000111100100011110010001111001000111100100011110000001111000000111100000011110000001110111000111011100011101110001110111000111011100011101100001110110000111011000011101010001110101000111010100011101010001110100000111010000011101000001110100000111001100011100110001110011000111001000011100100001110010000111000100011100010001110001000111000000011100000001110000000111000000011011110001101111000110111100011011100001101110000110111000011011010001101101000110110000011011000001101100000110101100011010110001101011000110101000011010100001101010000110100100011010010001101001000110100000011010000001100111000110011100011001110001100110000110011000011001010001100101000110010100011001000001100100000110001100011000110001100011000110001000011000100001100001000110000100011000010001100000000110000000010111110001011111000101111100010111100001011110000101110100010111010001011100000101110000010111000001011011000101101100010110100001011010000101100100010110010001011001000101100000010110000001010111000101011100010101100001010110000101010100010101010001010101000101010000010101000001010011000101001100010100100001010010000101000100010100010001010001000101000000010100000001001111000100111100010011100001001110000100110100010011010001001101000100110000010011000001001011000100101100010010100001001010000100100100010010010001001000000100100000010010000001000111000100011100010001100001000110000100010100010001010001000100000100010000010000110001000011000100001100010000100001000010000100000100010000010001000000000100000000001111110000111111000011111100001111100000111110000011110100001111010000111100000011110000001110110000111011000011101100001110100000111010000011100100001110010000111000000011100000001110000000110111000011011100001101100000110110000011010100001101010000110101000011010000001101000000110011000011001100001100100000110010000011001000001100010000110001000011000000001100000000110000000010111100001011110000101110000010111000001011100000101101000010110100001011000000101100000010110000001010110000101011000010101000001010100000101010000010100100001010010000101000000010100000001010000000100111000010011100001001110000100110000010011000001001010000100101000010010100001001000000100100000010010000001000110000100011000010001100001000100000100010000010000100001000010000100001000010000000001000000000100000000001111100000111110000011111000001111000000111100000011110000001110100000111010000011101000001110000000111000000011100000001101100000110110000011011000001101100000110100000011010000001101000000110010000011001000001100100000110000000011000000001100000000110000000010111000001011100000101110000010110000001011000000101100000010110000001010100000101010000010101000001010000000101000000010100000001010000000100110000010011000001001100000100110000010010000001001000000100100000010010000001000100000100010000010001000001000100000100000000010000000001000000000100000000010000000000111100000011110000001111000000111100000011100000001110000000111000000011100000001110000000110100000011010000001101000000110100000011010000001100000000110000000011000000001100000000110000000010110000001011000000101100000010110000001011000000101100000010100000001010000000101000000010100000001010000000100100000010010000001001000000100100000010010000001001000000100000000010000000001000000000100000000010000000001000000000100000000001110000000111000000011100000001110000000111000000011100000001110000000110000000011000000001100000000110000000011000000001100000000110000000011000000001010000000101000000010100000001010000000101000000010100000001010000000101000000010100000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111; 
        endcase      
    end
    else if (i_WIND_sel == NB_SEL'b11) begin // Kaiser with B = 14
        case (i_NFFT_sel)
            3'b000 : o_window = 160'b0000000000000000000000000000010000001000000001101100001110110001100001000111110000011111000001100001000011101100000110110000001000000000000100000000000000000000;
            3'b001 : o_window = 320'b00000000000000000000000000000000000000000000000001000000001100000001110000001110000001011100001001000000110101000100011100010110100001101011000111100000011111110001111111000111100000011010110001011010000100011100001101010000100100000001011100000011100000000111000000001100000000010000000000000000000000000000000000000000;
            3'b010 : o_window = 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000001100000001010000000111000000100100000011010000010001000001011000000111000000100010000010101000001100100000111011000100010000010011010001010110000101111100011010000001101111000111010100011110100001111110000111111100011111110001111110000111101000011101010001101111000110100000010111110001010110000100110100010001000000111011000011001000001010100000100010000001110000000101100000010001000000110100000010010000000111000000010100000000110000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
            3'b011 : o_window = 1280'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000100000000100000000010000000001100000001000000000100000000010100000001100000001000000000100100000010110000001100000000111000000100000000010011000001010100000110000000011011000001111000001000010000100101000010100100001011010000110001000011010100001110010000111110000100001000010001110001001011000101000000010101010001011001000101111000011000100001100110000110101000011011010001110001000111010000011101110001111001000111101100011111010001111110000111111100011111110001111111000111111100011111100001111101000111101100011110010001110111000111010000011100010001101101000110101000011001100001100010000101111000010110010001010101000101000000010010110001000111000100001000001111100000111001000011010100001100010000101101000010100100001001010000100001000001111000000110110000011000000001010100000100110000010000000000111000000011000000001011000000100100000010000000000110000000010100000001000000000100000000001100000000100000000010000000000100000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            3'b100 : o_window = 2560'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000010000000001000000000100000000010000000010000000001000000000100000000010000000001100000000110000000100000000010000000001000000000101000000010100000001100000000110000000011100000010000000001000000000100100000010100000001010000000101100000011000000001101000000111000000011110000010000000001000100000100100000010100000001010100000101100000011000000001100100000110110000011100000001111000000111110000100001000010001100001001000000100110000010100000001010100000101100000010111000001100000000110010000011010000001101100000111001000011101100001111010000111111000100000100010001000001000110000100100000010010110001001101000100111100010100010001010100000101011000010110000001011010000101110100010111110001100001000110001100011001010001100111000110100100011010110001101101000110111000011100000001110010000111001100011101010001110110000111011100011110010001111010000111101100011111000001111101000111110100011111100001111110000111111100011111110001111111000111111100011111110001111111000111111100011111110001111110000111111000011111010001111101000111110000011110110001111010000111100100011101110001110110000111010100011100110001110010000111000000011011100001101101000110101100011010010001100111000110010100011000110001100001000101111100010111010001011010000101100000010101100001010100000101000100010011110001001101000100101100010010000001000110000100010000010000010000111111000011110100001110110000111001000011011000001101000000110010000011000000001011100000101100000010101000001010000000100110000010010000001000110000100001000001111100000111100000011100000001101100000110010000011000000001011000000101010000010100000001001000000100010000010000000000111100000011100000001101000000110000000010110000001010000000101000000010010000001000000000100000000001110000000110000000011000000001010000000101000000010000000001000000000100000000001100000000110000000010000000001000000000100000000010000000000100000000010000000001000000000100000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            3'b101 : o_window = 5120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000001000000000100000000010000000001000000000100000000010000000001000000000100000000011000000001100000000110000000011000000001100000000110000000100000000010000000001000000000100000000010100000001010000000101000000010100000001010000000110000000011000000001100000000111000000011100000001110000000111000000100000000010000000001001000000100100000010010000001010000000101000000010100000001011000000101100000011000000001100000000110100000011010000001101000000111000000011100000001111000000111100000100000000010001000001000100000100100000010010000001001100000101000000010100000001010100000101010000010110000001011100000101110000011000000001100100000110100000011010000001101100000111000000011101000001110100000111100000011111000010000000001000010000100010000010001000001000110000100100000010010100001001100000100111000010100000001010010000101010000010101100001011000000101101000010111000001011110000110000000011000100001100100000110011000011010000001101010000110110000011011100001110000000111001000011101000001110110000111101000011111000001111110001000000000100000100010000100001000011000100010000010001100001000111000100100000010010010001001010000100101100010011000001001110000100111100010100000001010001000101001000010100110001010100000101011000010101110001011000000101100100010110100001011011000101110000010111010001011110000101111100011000010001100010000110001100011001000001100101000110011000011001110001101000000110100100011010100001101011000110101100011011000001101101000110111000011011110001110000000111000100011100010001110010000111001100011101000001110100000111010100011101100001110111000111011100011110000001111000000111100100011110100001111010000111101100011110110001111100000111110000011111000001111101000111110100011111010001111110000111111000011111100001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111110000111111000011111100001111101000111110100011111010001111100000111110000011111000001111011000111101100011110100001111010000111100100011110000001111000000111011100011101110001110110000111010100011101000001110100000111001100011100100001110001000111000100011100000001101111000110111000011011010001101100000110101100011010110001101010000110100100011010000001100111000110011000011001010001100100000110001100011000100001100001000101111100010111100001011101000101110000010110110001011010000101100100010110000001010111000101011000010101000001010011000101001000010100010001010000000100111100010011100001001100000100101100010010100001001001000100100000010001110001000110000100010000010000110001000010000100000100010000000000111111000011111000001111010000111011000011101000001110010000111000000011011100001101100000110101000011010000001100110000110010000011000100001100000000101111000010111000001011010000101100000010101100001010100000101001000010100000001001110000100110000010010100001001000000100011000010001000001000100000100001000010000000000111110000011110000001110100000111010000011100000001101100000110100000011010000001100100000110000000010111000001011100000101100000010101000001010100000101000000010100000001001100000100100000010010000001000100000100010000010000000000111100000011110000001110000000111000000011010000001101000000110100000011000000001100000000101100000010110000001010000000101000000010100000001001000000100100000010010000001000000000100000000001110000000111000000011100000001110000000110000000011000000001100000000101000000010100000001010000000101000000010100000001000000000100000000010000000001000000000011000000001100000000110000000011000000001100000000110000000010000000001000000000100000000010000000001000000000100000000010000000001000000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            3'b110 : o_window = 10240'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001010000000101000000010100000001010000000101000000010100000001010000000101000000011000000001100000000110000000011000000001100000000110000000011000000001110000000111000000011100000001110000000111000000011100000001110000001000000000100000000010000000001000000000100000000010000000001001000000100100000010010000001001000000100100000010100000001010000000101000000010100000001010000000101100000010110000001011000000101100000010110000001100000000110000000011000000001100000000110000000011010000001101000000110100000011010000001110000000111000000011100000001110000000111100000011110000001111000000111100000100000000010000000001000000000100010000010001000001000100000100010000010010000001001000000100100000010011000001001100000100110000010011000001010000000101000000010100000001010100000101010000010101000001011000000101100000010110000001011100000101110000010111000001100000000110000000011000000001100100000110010000011001000001101000000110100000011011000001101100000110110000011100000001110000000111010000011101000001110100000111100000011110000001111100000111110000011111000010000000001000000000100001000010000100001000010000100010000010001000001000110000100011000010010000001001000000100100000010010100001001010000100110000010011000001001110000100111000010100000001010000000101001000010100100001010100000101010000010101100001010110000101100000010110000001011010000101101000010111000001011100000101111000010111100001100000000110000000011000100001100010000110010000011001000001100110000110011000011010000001101000000110101000011010100001101100000110110000011011100001101110000111000000011100100001110010000111010000011101000001110110000111011000011110000001111000000111101000011111000001111100000111111000011111100010000000001000000000100000100010000010001000010000100001100010000110001000100000100010000010001010001000101000100011000010001110001000111000100100000010010000001001001000100100100010010100001001011000100101100010011000001001100000100110100010011010001001110000100111100010011110001010000000101000000010100010001010001000101001000010100110001010011000101010000010101000001010101000101010100010101100001010111000101011100010110000001011000000101100100010110010001011010000101101000010110110001011100000101110000010111010001011101000101111000010111100001011111000101111100011000000001100000000110000100011000010001100010000110001000011000110001100011000110010000011001000001100101000110010100011001100001100110000110011100011001110001101000000110100000011010010001101001000110101000011010100001101011000110101100011011000001101100000110110100011011010001101101000110111000011011100001101111000110111100011100000001110000000111000000011100010001110001000111001000011100100001110010000111001100011100110001110100000111010000011101000001110101000111010100011101010001110110000111011000011101100001110111000111011100011101110001111000000111100000011110000001111001000111100100011110010001111001000111101000011110100001111010000111101000011110110001111011000111101100011110110001111100000111110000011111000001111100000111110000011111010001111101000111110100011111010001111101000111111000011111100001111110000111111000011111100001111110000111111000011111100001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111100011111110001111111000111111000011111100001111110000111111000011111100001111110000111111000011111100001111101000111110100011111010001111101000111110100011111000001111100000111110000011111000001111100000111101100011110110001111011000111101100011110100001111010000111101000011110100001111001000111100100011110010001111001000111100000011110000001111000000111011100011101110001110111000111011000011101100001110110000111010100011101010001110101000111010000011101000001110100000111001100011100110001110010000111001000011100100001110001000111000100011100000001110000000111000000011011110001101111000110111000011011100001101101000110110100011011010001101100000110110000011010110001101011000110101000011010100001101001000110100100011010000001101000000110011100011001110001100110000110011000011001010001100101000110010000011001000001100011000110001100011000100001100010000110000100011000010001100000000110000000010111110001011111000101111000010111100001011101000101110100010111000001011100000101101100010110100001011010000101100100010110010001011000000101100000010101110001010111000101011000010101010001010101000101010000010101000001010011000101001100010100100001010001000101000100010100000001010000000100111100010011110001001110000100110100010011010001001100000100110000010010110001001011000100101000010010010001001001000100100000010010000001000111000100011100010001100001000101000100010100010001000001000100000100001100010000110001000010000100000100010000010001000000000100000000001111110000111111000011111000001111100000111101000011110000001111000000111011000011101100001110100000111010000011100100001110010000111000000011011100001101110000110110000011011000001101010000110101000011010000001101000000110011000011001100001100100000110010000011000100001100010000110000000011000000001011110000101111000010111000001011100000101101000010110100001011000000101100000010101100001010110000101010000010101000001010010000101001000010100000001010000000100111000010011100001001100000100110000010010100001001010000100100000010010000001001000000100011000010001100001000100000100010000010000100001000010000100001000010000000001000000000011111000001111100000111110000011110000001111000000111010000011101000001110100000111000000011100000001101100000110110000011011000001101000000110100000011001000001100100000110010000011000000001100000000110000000010111000001011100000101110000010110000001011000000101100000010101000001010100000101010000010100000001010000000101000000010011000001001100000100110000010011000001001000000100100000010010000001000100000100010000010001000001000100000100000000010000000001000000000011110000001111000000111100000011110000001110000000111000000011100000001110000000110100000011010000001101000000110100000011000000001100000000110000000011000000001100000000101100000010110000001011000000101100000010110000001010000000101000000010100000001010000000101000000010010000001001000000100100000010010000001001000000100000000010000000001000000000100000000010000000001000000000011100000001110000000111000000011100000001110000000111000000011100000001100000000110000000011000000001100000000110000000011000000001100000000101000000010100000001010000000101000000010100000001010000000101000000010100000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; 
        endcase       
    end  
end

endmodule